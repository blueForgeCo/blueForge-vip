
package base_test_lib_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "components/base_env.svh"
    `include "components/base_component.svh"

endpackage

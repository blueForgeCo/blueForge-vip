
package bforge_apb_lib_pkg;

    import uvm_pkg::*;
    import bforge_base_lib_pkg::*;
    `include "uvm_macros.svh"

    `include "types/apb_types.svh"
    `include "types/apb_config.svh"

    `include "seq_items/apb_txn.svh"

    `include "components/apb_sequencer.svh"
    `include "components/apb_driver.svh"
    `include "components/apb_monitor.svh"
    `include "components/apb_agent.svh"

endpackage

`include "interfaces/bforge_apb_if.sv"
`include "modules/bforge_apb_initiator.sv"
`include "modules/bforge_apb_monitor.sv"
`include "modules/bforge_apb_target.sv"


package params_pkg;

    parameter int TARGET_COUNT = 4;

endpackage


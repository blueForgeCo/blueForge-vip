
package params_pkg;

    parameter int TARGET_COUNT = 5;

endpackage


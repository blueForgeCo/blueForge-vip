
package bforge_base_lib_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "types/base_types.svh"
    `include "components/base_agent.svh"
    `include "components/base_driver.svh"
    `include "components/base_monitor.svh"

endpackage

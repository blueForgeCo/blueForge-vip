
typedef bit[63:00] addr_t;
typedef bit[04:00] int4_t;
typedef bit[07:00] int8_t;
typedef bit[16:00] int16_t;
typedef bit[31:00] int32_t;
typedef bit[63:00] int64_t;

